-------------------------------------------------------------------------------
--
-- Title       : No Title
-- Design      : projeto06281
-- Author      : julia.fernandes.moraes@usp.br
-- Company     : usp
--
-------------------------------------------------------------------------------
--
-- File        : C:\My_Designs\projeto1\projeto06281\compile\uc+hierarquia.vhd
-- Generated   : Sun Jun 30 20:11:39 2019
-- From        : C:/My_Designs/projeto1/projeto06281/src/uc+hierarquia.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_unsigned.all;

entity \uc+hierarquia\ is 
end \uc+hierarquia\;

architecture \uc+hierarquia\ of \uc+hierarquia\ is

---- Component declarations -----

component Fub1
	--- component Fub1 has no ports
end component;
component Fub2
	--- component Fub2 has no ports
end component;

begin

----  Component instantiations  ----

U1 : Fub1;

U2 : Fub2;


end \uc+hierarquia\;
